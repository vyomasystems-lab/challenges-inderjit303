
module PGGen(output g, p, input a, b);
 
  and #(1) (g, a, b);
  xor #(2) (p, a, b);
 
endmodule

module CLA32(output [31:0] sum, output cout, input [31:0] a, b);
wire [31:0] g, p, c;
wire [1000:0] e;
wire cin;
buf #(1) (cin, 0);
//c[0]
and #(1) (e[0], cin, p[0]);
or #(1) (c[0], e[0], g[0]);

//c[1]
and #(1) (e[1], cin, p[0], p[1]);
and #(1) (e[2], g[0], p[1]);
or #(1) (c[1], e[1], e[2], g[1]);

//c[2]
and #(1) (e[3], cin, p[0], p[1], p[2]);
and #(1) (e[4], g[0], p[1], p[2]);
and #(1) (e[5], g[1], p[2]);
or #(1) (c[2], e[3], e[4], e[5], g[2]);

//c[3]
and #(1) (e[6], cin, p[0], p[1], p[2], p[3]);
and #(1) (e[7], g[0], p[1], p[2], p[3]);
and #(1) (e[8], g[1], p[2], p[3]);
and #(1) (e[9], g[2], p[3]);
or #(1) (c[3], e[6], e[7], e[8], e[9], g[3]);

//c[4]
and #(1) (e[10], cin, p[0], p[1], p[2], p[3], p[4]);
and #(1) (e[11], g[0], p[1], p[2], p[3], p[4]);
and #(1) (e[12], g[1], p[2], p[3], p[4]);
and #(1) (e[13], g[2], p[3], p[4]);
and #(1) (e[14], g[3], p[4]);
or #(1) (c[4], e[10], e[11], e[12], e[13], e[14], g[4]);

//c[5]
and #(1) (e[15], cin, p[0], p[1], p[2], p[3], p[4], p[5]);
and #(1) (e[16], g[0], p[1], p[2], p[3], p[4], p[5]);
and #(1) (e[17], g[1], p[2], p[3], p[4], p[5]);
and #(1) (e[18], g[2], p[3], p[4], p[5]);
and #(1) (e[19], g[3], p[4], p[5]);
and #(1) (e[20], g[4], p[5]);
or #(1) (c[5], e[15], e[16], e[17], e[18], e[19], e[20], g[5]);

//c[6]
and #(1) (e[21], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6]);
and #(1) (e[22], g[0], p[1], p[2], p[3], p[4], p[5], p[6]);
and #(1) (e[23], g[1], p[2], p[3], p[4], p[5], p[6]);
and #(1) (e[24], g[2], p[3], p[4], p[5], p[6]);
and #(1) (e[25], g[3], p[4], p[5], p[6]);
and #(1) (e[26], g[4], p[5], p[6]);
and #(1) (e[27], g[5], p[6]);
or #(1) (c[6], e[21], e[22], e[23], e[24], e[25], e[26], e[27], g[6]);

//c[7]
and #(1) (e[28], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7]);
and #(1) (e[29], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7]);
and #(1) (e[30], g[1], p[2], p[3], p[4], p[5], p[6], p[7]);
and #(1) (e[31], g[2], p[3], p[4], p[5], p[6], p[7]);
and #(1) (e[32], g[3], p[4], p[5], p[6], p[7]);
and #(1) (e[33], g[4], p[5], p[6], p[7]);
and #(1) (e[34], g[5], p[6], p[7]);
and #(1) (e[35], g[6], p[7]);
or #(1) (c[7], e[28], e[29], e[30], e[31], e[32], e[33], e[34], e[35], g[7]);

//c[8]
and #(1) (e[36], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8]);
and #(1) (e[37], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8]);
and #(1) (e[38], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8]);
and #(1) (e[39], g[2], p[3], p[4], p[5], p[6], p[7], p[8]);
and #(1) (e[40], g[3], p[4], p[5], p[6], p[7], p[8]);
and #(1) (e[41], g[4], p[5], p[6], p[7], p[8]);
and #(1) (e[42], g[5], p[6], p[7], p[8]);
and #(1) (e[43], g[6], p[7], p[8]);
and #(1) (e[44], g[7], p[8]);
or #(1) (c[8], e[36], e[37], e[38], e[39], e[40], e[41], e[42], e[43], e[44], g[8]);

//c[9]
and #(1) (e[45], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9]);
and #(1) (e[46], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9]);
and #(1) (e[47], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9]);
and #(1) (e[48], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9]);
and #(1) (e[49], g[3], p[4], p[5], p[6], p[7], p[8], p[9]);
and #(1) (e[50], g[4], p[5], p[6], p[7], p[8], p[9]);
and #(1) (e[51], g[5], p[6], p[7], p[8], p[9]);
and #(1) (e[52], g[6], p[7], p[8], p[9]);
and #(1) (e[53], g[7], p[8], p[9]);
and #(1) (e[54], g[8], p[9]);
or #(1) (c[9], e[45], e[46], e[47], e[48], e[49], e[50], e[51], e[52], e[53], e[54], g[9]);

//c[10]
and #(1) (e[55], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10]);
and #(1) (e[56], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10]);
and #(1) (e[57], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10]);
and #(1) (e[58], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10]);
and #(1) (e[59], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10]);
and #(1) (e[60], g[4], p[5], p[6], p[7], p[8], p[9], p[10]);
and #(1) (e[61], g[5], p[6], p[7], p[8], p[9], p[10]);
and #(1) (e[62], g[6], p[7], p[8], p[9], p[10]);
and #(1) (e[63], g[7], p[8], p[9], p[10]);
and #(1) (e[64], g[8], p[9], p[10]);
and #(1) (e[65], g[9], p[10]);
or #(1) (c[10], e[55], e[56], e[57], e[58], e[59], e[60], e[61], e[62], e[63], e[64], e[65], g[10]);

//c[11]
and #(1) (e[66], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11]);
and #(1) (e[67], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11]);
and #(1) (e[68], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11]);
and #(1) (e[69], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11]);
and #(1) (e[70], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11]);
and #(1) (e[71], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11]);
and #(1) (e[72], g[5], p[6], p[7], p[8], p[9], p[10], p[11]);
and #(1) (e[73], g[6], p[7], p[8], p[9], p[10], p[11]);
and #(1) (e[74], g[7], p[8], p[9], p[10], p[11]);
and #(1) (e[75], g[8], p[9], p[10], p[11]);
and #(1) (e[76], g[9], p[10], p[11]);
and #(1) (e[77], g[10], p[11]);
or #(1) (c[11], e[66], e[67], e[68], e[69], e[70], e[71], e[72], e[73], e[74], e[75], e[76], e[77], g[11]);

//c[12]
and #(1) (e[78], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12]);
and #(1) (e[79], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12]);
and #(1) (e[80], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12]);
and #(1) (e[81], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12]);
and #(1) (e[82], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12]);
and #(1) (e[83], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12]);
and #(1) (e[84], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12]);
and #(1) (e[85], g[6], p[7], p[8], p[9], p[10], p[11], p[12]);
and #(1) (e[86], g[7], p[8], p[9], p[10], p[11], p[12]);
and #(1) (e[87], g[8], p[9], p[10], p[11], p[12]);
and #(1) (e[88], g[9], p[10], p[11], p[12]);
and #(1) (e[89], g[10], p[11], p[12]);
and #(1) (e[90], g[11], p[12]);
or #(1) (c[12], e[78], e[79], e[80], e[81], e[82], e[83], e[84], e[85], e[86], e[87], e[88], e[89], e[90], g[12]);

//c[13]
and #(1) (e[91], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13]);
and #(1) (e[92], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13]);
and #(1) (e[93], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13]);
and #(1) (e[94], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13]);
and #(1) (e[95], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13]);
and #(1) (e[96], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13]);
and #(1) (e[97], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13]);
and #(1) (e[98], g[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13]);
and #(1) (e[99], g[7], p[8], p[9], p[10], p[11], p[12], p[13]);
and #(1) (e[100], g[8], p[9], p[10], p[11], p[12], p[13]);
and #(1) (e[101], g[9], p[10], p[11], p[12], p[13]);
and #(1) (e[102], g[10], p[11], p[12], p[13]);
and #(1) (e[103], g[11], p[12], p[13]);
and #(1) (e[104], g[12], p[13]);
or #(1) (c[13], e[91], e[92], e[93], e[94], e[95], e[96], e[97], e[98], e[99], e[100], e[101], e[102], e[103], e[104], g[13]);

//c[14]
and #(1) (e[105], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14]);
and #(1) (e[106], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14]);
and #(1) (e[107], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14]);
and #(1) (e[108], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14]);
and #(1) (e[109], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14]);
and #(1) (e[110], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14]);
and #(1) (e[111], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14]);
and #(1) (e[112], g[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14]);
and #(1) (e[113], g[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14]);
and #(1) (e[114], g[8], p[9], p[10], p[11], p[12], p[13], p[14]);
and #(1) (e[115], g[9], p[10], p[11], p[12], p[13], p[14]);
and #(1) (e[116], g[10], p[11], p[12], p[13], p[14]);
and #(1) (e[117], g[11], p[12], p[13], p[14]);
and #(1) (e[118], g[12], p[13], p[14]);
and #(1) (e[119], g[13], p[14]);
or #(1) (c[14], e[105], e[106], e[107], e[108], e[109], e[110], e[111], e[112], e[113], e[114], e[115], e[116], e[117], e[118], e[119], g[14]);

//c[15]
and #(1) (e[120], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[121], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[122], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[123], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[124], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[125], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[126], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[127], g[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[128], g[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[129], g[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[130], g[9], p[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[131], g[10], p[11], p[12], p[13], p[14], p[15]);
and #(1) (e[132], g[11], p[12], p[13], p[14], p[15]);
and #(1) (e[133], g[12], p[13], p[14], p[15]);
and #(1) (e[134], g[13], p[14], p[15]);
and #(1) (e[135], g[14], p[15]);
or #(1) (c[15], e[120], e[121], e[122], e[123], e[124], e[125], e[126], e[127], e[128], e[129], e[130], e[131], e[132], e[133], e[134], e[135], g[15]);

//c[16]
and #(1) (e[136], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16]);
and #(1) (e[137], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16]);
and #(1) (e[138], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16]);
and #(1) (e[139], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16]);
and #(1) (e[140], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16]);
and #(1) (e[141], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16]);
and #(1) (e[142], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16]);
and #(1) (e[143], g[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16]);
and #(1) (e[144], g[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16]);
and #(1) (e[145], g[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16]);
and #(1) (e[146], g[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16]);
and #(1) (e[147], g[10], p[11], p[12], p[13], p[14], p[15], p[16]);
and #(1) (e[148], g[11], p[12], p[13], p[14], p[15], p[16]);
and #(1) (e[149], g[12], p[13], p[14], p[15], p[16]);
and #(1) (e[150], g[13], p[14], p[15], p[16]);
and #(1) (e[151], g[14], p[15], p[16]);
and #(1) (e[152], g[15], p[16]);
or #(1) (c[16], e[136], e[137], e[138], e[139], e[140], e[141], e[142], e[143], e[144], e[145], e[146], e[147], e[148], e[149], e[150], e[151], e[152], g[16]);

//c[17]
and #(1) (e[153], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17]);
and #(1) (e[154], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17]);
and #(1) (e[155], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17]);
and #(1) (e[156], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17]);
and #(1) (e[157], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17]);
and #(1) (e[158], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17]);
and #(1) (e[159], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17]);
and #(1) (e[160], g[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17]);
and #(1) (e[161], g[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17]);
and #(1) (e[162], g[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17]);
and #(1) (e[163], g[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17]);
and #(1) (e[164], g[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17]);
and #(1) (e[165], g[11], p[12], p[13], p[14], p[15], p[16], p[17]);
and #(1) (e[166], g[12], p[13], p[14], p[15], p[16], p[17]);
and #(1) (e[167], g[13], p[14], p[15], p[16], p[17]);
and #(1) (e[168], g[14], p[15], p[16], p[17]);
and #(1) (e[169], g[15], p[16], p[17]);
and #(1) (e[170], g[16], p[17]);
or #(1) (c[17], e[153], e[154], e[155], e[156], e[157], e[158], e[159], e[160], e[161], e[162], e[163], e[164], e[165], e[166], e[167], e[168], e[169], e[170], g[17]);

//c[18]
and #(1) (e[171], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18]);
and #(1) (e[172], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18]);
and #(1) (e[173], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18]);
and #(1) (e[174], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18]);
and #(1) (e[175], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18]);
and #(1) (e[176], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18]);
and #(1) (e[177], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18]);
and #(1) (e[178], g[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18]);
and #(1) (e[179], g[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18]);
and #(1) (e[180], g[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18]);
and #(1) (e[181], g[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18]);
and #(1) (e[182], g[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18]);
and #(1) (e[183], g[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18]);
and #(1) (e[184], g[12], p[13], p[14], p[15], p[16], p[17], p[18]);
and #(1) (e[185], g[13], p[14], p[15], p[16], p[17], p[18]);
and #(1) (e[186], g[14], p[15], p[16], p[17], p[18]);
and #(1) (e[187], g[15], p[16], p[17], p[18]);
and #(1) (e[188], g[16], p[17], p[18]);
and #(1) (e[189], g[17], p[18]);
or #(1) (c[18], e[171], e[172], e[173], e[174], e[175], e[176], e[177], e[178], e[179], e[180], e[181], e[182], e[183], e[184], e[185], e[186], e[187], e[188], e[189], g[18]);

//c[19]
and #(1) (e[190], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19]);
and #(1) (e[191], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19]);
and #(1) (e[192], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19]);
and #(1) (e[193], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19]);
and #(1) (e[194], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19]);
and #(1) (e[195], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19]);
and #(1) (e[196], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19]);
and #(1) (e[197], g[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19]);
and #(1) (e[198], g[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19]);
and #(1) (e[199], g[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19]);
and #(1) (e[200], g[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19]);
and #(1) (e[201], g[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19]);
and #(1) (e[202], g[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19]);
and #(1) (e[203], g[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19]);
and #(1) (e[204], g[13], p[14], p[15], p[16], p[17], p[18], p[19]);
and #(1) (e[205], g[14], p[15], p[16], p[17], p[18], p[19]);
and #(1) (e[206], g[15], p[16], p[17], p[18], p[19]);
and #(1) (e[207], g[16], p[17], p[18], p[19]);
and #(1) (e[208], g[17], p[18], p[19]);
and #(1) (e[209], g[18], p[19]);
or #(1) (c[19], e[190], e[191], e[192], e[193], e[194], e[195], e[196], e[197], e[198], e[199], e[200], e[201], e[202], e[203], e[204], e[205], e[206], e[207], e[208], e[209], g[19]);

//c[20]
and #(1) (e[210], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20]);
and #(1) (e[211], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20]);
and #(1) (e[212], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20]);
and #(1) (e[213], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20]);
and #(1) (e[214], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20]);
and #(1) (e[215], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20]);
and #(1) (e[216], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20]);
and #(1) (e[217], g[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20]);
and #(1) (e[218], g[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20]);
and #(1) (e[219], g[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20]);
and #(1) (e[220], g[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20]);
and #(1) (e[221], g[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20]);
and #(1) (e[222], g[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20]);
and #(1) (e[223], g[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20]);
and #(1) (e[224], g[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20]);
and #(1) (e[225], g[14], p[15], p[16], p[17], p[18], p[19], p[20]);
and #(1) (e[226], g[15], p[16], p[17], p[18], p[19], p[20]);
and #(1) (e[227], g[16], p[17], p[18], p[19], p[20]);
and #(1) (e[228], g[17], p[18], p[19], p[20]);
and #(1) (e[229], g[18], p[19], p[20]);
and #(1) (e[230], g[19], p[20]);
or #(1) (c[20], e[210], e[211], e[212], e[213], e[214], e[215], e[216], e[217], e[218], e[219], e[220], e[221], e[222], e[223], e[224], e[225], e[226], e[227], e[228], e[229], e[230], g[20]);

//c[21]
and #(1) (e[231], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21]);
and #(1) (e[232], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21]);
and #(1) (e[233], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21]);
and #(1) (e[234], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21]);
and #(1) (e[235], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21]);
and #(1) (e[236], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21]);
and #(1) (e[237], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21]);
and #(1) (e[238], g[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21]);
and #(1) (e[239], g[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21]);
and #(1) (e[240], g[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21]);
and #(1) (e[241], g[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21]);
and #(1) (e[242], g[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21]);
and #(1) (e[243], g[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21]);
and #(1) (e[244], g[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21]);
and #(1) (e[245], g[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21]);
and #(1) (e[246], g[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21]);
and #(1) (e[247], g[15], p[16], p[17], p[18], p[19], p[20], p[21]);
and #(1) (e[248], g[16], p[17], p[18], p[19], p[20], p[21]);
and #(1) (e[249], g[17], p[18], p[19], p[20], p[21]);
and #(1) (e[250], g[18], p[19], p[20], p[21]);
and #(1) (e[251], g[19], p[20], p[21]);
and #(1) (e[252], g[20], p[21]);
or #(1) (c[21], e[231], e[232], e[233], e[234], e[235], e[236], e[237], e[238], e[239], e[240], e[241], e[242], e[243], e[244], e[245], e[246], e[247], e[248], e[249], e[250], e[251], e[252], g[21]);

//c[22]
and #(1) (e[253], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22]);
and #(1) (e[254], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22]);
and #(1) (e[255], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22]);
and #(1) (e[256], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22]);
and #(1) (e[257], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22]);
and #(1) (e[258], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22]);
and #(1) (e[259], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22]);
and #(1) (e[260], g[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22]);
and #(1) (e[261], g[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22]);
and #(1) (e[262], g[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22]);
and #(1) (e[263], g[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22]);
and #(1) (e[264], g[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22]);
and #(1) (e[265], g[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22]);
and #(1) (e[266], g[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22]);
and #(1) (e[267], g[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22]);
and #(1) (e[268], g[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22]);
and #(1) (e[269], g[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22]);
and #(1) (e[270], g[16], p[17], p[18], p[19], p[20], p[21], p[22]);
and #(1) (e[271], g[17], p[18], p[19], p[20], p[21], p[22]);
and #(1) (e[272], g[18], p[19], p[20], p[21], p[22]);
and #(1) (e[273], g[19], p[20], p[21], p[22]);
and #(1) (e[274], g[20], p[21], p[22]);
and #(1) (e[275], g[21], p[22]);
or #(1) (c[22], e[253], e[254], e[255], e[256], e[257], e[258], e[259], e[260], e[261], e[262], e[263], e[264], e[265], e[266], e[267], e[268], e[269], e[270], e[271], e[272], e[273], e[274], e[275], g[22]);

//c[23]
and #(1) (e[276], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23]);
and #(1) (e[277], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23]);
and #(1) (e[278], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23]);
and #(1) (e[279], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23]);
and #(1) (e[280], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23]);
and #(1) (e[281], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23]);
and #(1) (e[282], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23]);
and #(1) (e[283], g[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23]);
and #(1) (e[284], g[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23]);
and #(1) (e[285], g[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23]);
and #(1) (e[286], g[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23]);
and #(1) (e[287], g[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23]);
and #(1) (e[288], g[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23]);
and #(1) (e[289], g[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23]);
and #(1) (e[290], g[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23]);
and #(1) (e[291], g[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23]);
and #(1) (e[292], g[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23]);
and #(1) (e[293], g[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23]);
and #(1) (e[294], g[17], p[18], p[19], p[20], p[21], p[22], p[23]);
and #(1) (e[295], g[18], p[19], p[20], p[21], p[22], p[23]);
and #(1) (e[296], g[19], p[20], p[21], p[22], p[23]);
and #(1) (e[297], g[20], p[21], p[22], p[23]);
and #(1) (e[298], g[21], p[22], p[23]);
and #(1) (e[299], g[22], p[23]);
or #(1) (c[23], e[276], e[277], e[278], e[279], e[280], e[281], e[282], e[283], e[284], e[285], e[286], e[287], e[288], e[289], e[290], e[291], e[292], e[293], e[294], e[295], e[296], e[297], e[298], e[299], g[23]);

//c[24]
and #(1) (e[300], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24]);
and #(1) (e[301], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24]);
and #(1) (e[302], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24]);
and #(1) (e[303], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24]);
and #(1) (e[304], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24]);
and #(1) (e[305], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24]);
and #(1) (e[306], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24]);
and #(1) (e[307], g[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24]);
and #(1) (e[308], g[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24]);
and #(1) (e[309], g[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24]);
and #(1) (e[310], g[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24]);
and #(1) (e[311], g[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24]);
and #(1) (e[312], g[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24]);
and #(1) (e[313], g[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24]);
and #(1) (e[314], g[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24]);
and #(1) (e[315], g[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24]);
and #(1) (e[316], g[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24]);
and #(1) (e[317], g[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24]);
and #(1) (e[318], g[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24]);
and #(1) (e[319], g[18], p[19], p[20], p[21], p[22], p[23], p[24]);
and #(1) (e[320], g[19], p[20], p[21], p[22], p[23], p[24]);
and #(1) (e[321], g[20], p[21], p[22], p[23], p[24]);
and #(1) (e[322], g[21], p[22], p[23], p[24]);
and #(1) (e[323], g[22], p[23], p[24]);
and #(1) (e[324], g[23], p[24]);
or #(1) (c[24], e[300], e[301], e[302], e[303], e[304], e[305], e[306], e[307], e[308], e[309], e[310], e[311], e[312], e[313], e[314], e[315], e[316], e[317], e[318], e[319], e[320], e[321], e[322], e[323], e[324], g[24]);

//c[25]
and #(1) (e[325], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25]);
and #(1) (e[326], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25]);
and #(1) (e[327], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25]);
and #(1) (e[328], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25]);
and #(1) (e[329], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25]);
and #(1) (e[330], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25]);
and #(1) (e[331], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25]);
and #(1) (e[332], g[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25]);
and #(1) (e[333], g[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25]);
and #(1) (e[334], g[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25]);
and #(1) (e[335], g[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25]);
and #(1) (e[336], g[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25]);
and #(1) (e[337], g[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25]);
and #(1) (e[338], g[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25]);
and #(1) (e[339], g[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25]);
and #(1) (e[340], g[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25]);
and #(1) (e[341], g[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25]);
and #(1) (e[342], g[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25]);
and #(1) (e[343], g[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25]);
and #(1) (e[344], g[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25]);
and #(1) (e[345], g[19], p[20], p[21], p[22], p[23], p[24], p[25]);
and #(1) (e[346], g[20], p[21], p[22], p[23], p[24], p[25]);
and #(1) (e[347], g[21], p[22], p[23], p[24], p[25]);
and #(1) (e[348], g[22], p[23], p[24], p[25]);
and #(1) (e[349], g[23], p[24], p[25]);
and #(1) (e[350], g[24], p[25]);
or #(1) (c[25], e[325], e[326], e[327], e[328], e[329], e[330], e[331], e[332], e[333], e[334], e[335], e[336], e[337], e[338], e[339], e[340], e[341], e[342], e[343], e[344], e[345], e[346], e[347], e[348], e[349], e[350], g[25]);

//c[26]
and #(1) (e[351], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26]);
and #(1) (e[352], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26]);
and #(1) (e[353], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26]);
and #(1) (e[354], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26]);
and #(1) (e[355], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26]);
and #(1) (e[356], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26]);
and #(1) (e[357], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26]);
and #(1) (e[358], g[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26]);
and #(1) (e[359], g[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26]);
and #(1) (e[360], g[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26]);
and #(1) (e[361], g[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26]);
and #(1) (e[362], g[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26]);
and #(1) (e[363], g[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26]);
and #(1) (e[364], g[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26]);
and #(1) (e[365], g[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26]);
and #(1) (e[366], g[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26]);
and #(1) (e[367], g[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26]);
and #(1) (e[368], g[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26]);
and #(1) (e[369], g[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26]);
and #(1) (e[370], g[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26]);
and #(1) (e[371], g[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26]);
and #(1) (e[372], g[20], p[21], p[22], p[23], p[24], p[25], p[26]);
and #(1) (e[373], g[21], p[22], p[23], p[24], p[25], p[26]);
and #(1) (e[374], g[22], p[23], p[24], p[25], p[26]);
and #(1) (e[375], g[23], p[24], p[25], p[26]);
and #(1) (e[376], g[24], p[25], p[26]);
and #(1) (e[377], g[25], p[26]);
or #(1) (c[26], e[351], e[352], e[353], e[354], e[355], e[356], e[357], e[358], e[359], e[360], e[361], e[362], e[363], e[364], e[365], e[366], e[367], e[368], e[369], e[370], e[371], e[372], e[373], e[374], e[375], e[376], e[377], g[26]);

//c[27]
and #(1) (e[378], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[379], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[380], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[381], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[382], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[383], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[384], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[385], g[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[386], g[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[387], g[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[388], g[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[389], g[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[390], g[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[391], g[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[392], g[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[393], g[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[394], g[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[395], g[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[396], g[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[397], g[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[398], g[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[399], g[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[400], g[21], p[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[401], g[22], p[23], p[24], p[25], p[26], p[27]);
and #(1) (e[402], g[23], p[24], p[25], p[26], p[27]);
and #(1) (e[403], g[24], p[25], p[26], p[27]);
and #(1) (e[404], g[25], p[26], p[27]);
and #(1) (e[405], g[26], p[27]);
or #(1) (c[27], e[378], e[379], e[380], e[381], e[382], e[383], e[384], e[385], e[386], e[387], e[388], e[389], e[390], e[391], e[392], e[393], e[394], e[395], e[396], e[397], e[398], e[399], e[400], e[401], e[402], e[403], e[404], e[405], g[27]);

//c[28]
and #(1) (e[406], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[407], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[408], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[409], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[410], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[411], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[412], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[413], g[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[414], g[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[415], g[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[416], g[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[417], g[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[418], g[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[419], g[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[420], g[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[421], g[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[422], g[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[423], g[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[424], g[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[425], g[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[426], g[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[427], g[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[428], g[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[429], g[22], p[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[430], g[23], p[24], p[25], p[26], p[27], p[28]);
and #(1) (e[431], g[24], p[25], p[26], p[27], p[28]);
and #(1) (e[432], g[25], p[26], p[27], p[28]);
and #(1) (e[433], g[26], p[27], p[28]);
and #(1) (e[434], g[27], p[28]);
or #(1) (c[28], e[406], e[407], e[408], e[409], e[410], e[411], e[412], e[413], e[414], e[415], e[416], e[417], e[418], e[419], e[420], e[421], e[422], e[423], e[424], e[425], e[426], e[427], e[428], e[429], e[430], e[431], e[432], e[433], e[434], g[28]);

//c[29]
and #(1) (e[435], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[436], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[437], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[438], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[439], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[440], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[441], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[442], g[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[443], g[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[444], g[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[445], g[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[446], g[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[447], g[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[448], g[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[449], g[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[450], g[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[451], g[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[452], g[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[453], g[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[454], g[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[455], g[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[456], g[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[457], g[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[458], g[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[459], g[23], p[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[460], g[24], p[25], p[26], p[27], p[28], p[29]);
and #(1) (e[461], g[25], p[26], p[27], p[28], p[29]);
and #(1) (e[462], g[26], p[27], p[28], p[29]);
and #(1) (e[463], g[27], p[28], p[29]);
and #(1) (e[464], g[28], p[29]);
or #(1) (c[29], e[435], e[436], e[437], e[438], e[439], e[440], e[441], e[442], e[443], e[444], e[445], e[446], e[447], e[448], e[449], e[450], e[451], e[452], e[453], e[454], e[455], e[456], e[457], e[458], e[459], e[460], e[461], e[462], e[463], e[464], g[29]);

//c[30]
and #(1) (e[465], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[466], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[467], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[468], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[469], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[470], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[471], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[472], g[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[473], g[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[474], g[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[475], g[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[476], g[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[477], g[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[478], g[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[479], g[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[480], g[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[481], g[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[482], g[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[483], g[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[484], g[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[485], g[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[486], g[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[487], g[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[488], g[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[489], g[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[490], g[24], p[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[491], g[25], p[26], p[27], p[28], p[29], p[30]);
and #(1) (e[492], g[26], p[27], p[28], p[29], p[30]);
and #(1) (e[493], g[27], p[28], p[29], p[30]);
and #(1) (e[494], g[28], p[29], p[30]);
and #(1) (e[495], g[29], p[30]);
or #(1) (c[30], e[465], e[466], e[467], e[468], e[469], e[470], e[471], e[472], e[473], e[474], e[475], e[476], e[477], e[478], e[479], e[480], e[481], e[482], e[483], e[484], e[485], e[486], e[487], e[488], e[489], e[490], e[491], e[492], e[493], e[494], e[495], g[30]);

//c[31]
and #(1) (e[496], cin, p[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[497], g[0], p[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[498], g[1], p[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[499], g[2], p[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[500], g[3], p[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[501], g[4], p[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[502], g[5], p[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[503], g[6], p[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[504], g[7], p[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[505], g[8], p[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[506], g[9], p[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[507], g[10], p[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[508], g[11], p[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[509], g[12], p[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[510], g[13], p[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[511], g[14], p[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[512], g[15], p[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[513], g[16], p[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[514], g[17], p[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[515], g[18], p[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[516], g[19], p[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[517], g[20], p[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[518], g[21], p[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[519], g[22], p[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[520], g[23], p[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[521], g[24], p[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[522], g[25], p[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[523], g[26], p[27], p[28], p[29], p[30], p[31]);
and #(1) (e[524], g[27], p[28], p[29], p[30], p[31]);
and #(1) (e[525], g[28], p[29], p[30], p[31]);
and #(1) (e[526], g[29], p[30], p[31]);
and #(1) (e[527], g[30], p[31]);
or #(1) (c[31], e[496], e[497], e[498], e[499], e[500], e[501], e[502], e[503], e[504], e[505], e[506], e[507], e[508], e[509], e[510], e[511], e[512], e[513], e[514], e[515], e[516], e[517], e[518], e[519], e[520], e[521], e[522], e[523], e[524], e[525], e[526], e[527], g[31]);

xor #(2) (sum[0],p[0],cin);
xor #(2) x[31:1](sum[31:1],p[31:1],c[30:0]);
buf #(1) (cout, c[31]);
PGGen pggen[31:0](g[31:0],p[31:0],a[31:0],b[31:0]);

endmodule
